module ex4(clock,X,Clear,C_32,C_31,C_30,C_29,C_28,C_27,C_26,C_25,C_24,C_23,C_22,C_21,C_20,C_19,C_18,C_17,C_16,C_15,C_14,C_13,C_12,C_11,C_10,C_9,C_8,C_7,C_6,C_5,C_4,C_3,C_2,C_1,C_0,W,Z);
input clock;
input X,Clear,C_32,C_31,C_30,C_29,C_28,C_27,C_26,C_25,C_24,C_23,C_22,C_21,C_20,C_19,C_18,C_17,C_16,C_15,C_14,C_13,C_12,C_11,C_10,C_9,C_8,C_7,C_6,C_5,C_4,C_3,C_2,C_1,C_0;
output W,Z;
reg S3,S2,S1,S0,S7,S6,S5,S4,S11,S10,S9,S8,S15,S14,S13,S12,S19,S18,S17,S16,S23,S22,S21,S20,S27,S26,S25,S24,S31,S30,S29,S28;
wire n134,n135,n136_1,n137,n138,n139,n140,n141_1,n142,n143,n144,n145,n146_1,n147,n148,n149,n150,n151_1,n152,n153,n154,n155,n156_1,n157,n158,n159,n160,n161_1,n162,n163,n164,n165,n166_1,n167,n168,n169,n170,n172,n173,n174,n175,n176_1,n177,n178,n179,n180,n181_1,n182,n183,n184,n185,n186_1,n187,n188,n189,n190,n191_1,n192,n193,n194,n195,n196_1,n197,n198,n199,n200,n201_1,n202,n203,n204,n205,n206_1,n207,n208,n209,n210,n211_1,n212,n213,n214,n215,n216_1,n217,n218,n219,n220,n221_1,n222,n223,n224,n225,n226_1,n227,n228,n229,n230,n231_1,n232,n233,n234,n235,n236,n237,n238,n239,n240,n241,n242,n243,n244,n245,n246,n247,n248,n249,n250,n251,n252,n253,n254,n255,n256,n257,n258,n259,n260,n261,n262,n263,n264,n265,n266,n267,n268,n269,n270,n271,n272,n273,n274,n275,n276,n277,n278,n279,n280,n281,n282,n283,n284,n285,n286,n287,n288,n289,n290,n291,n292,n293,n294,n295,n296,n297,n298,n299,n300,n301,n302,n303,n304,n305,n306,n307,n308,n309,n310,n311,n312,n313,n314,n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,n325,n326,n327,n328,n329,n330,n331,n332,n334,n335,n336,n337,n338,n339,n340,n341,n342,n343,n344,n345,n346,n347,n349,n350,n351,n352,n353,n354,n357,n358,n359,n360,n361,n363,n364,n365,n366,n367,n368,n369,n370,n371,n372,n373,n374,n375,n376,n377,n379,n380,n381,n382,n383,n384,n387,n388,n389,n390,n391,n393,n394,n395,n396,n397,n398,n399,n400,n401,n402,n403,n404,n405,n406,n407,n409,n410,n411,n412,n413,n414,n417,n418,n419,n420,n421,n423,n424,n425,n426,n427,n428,n429,n430,n431,n432,n433,n434,n435,n436,n437,n439,n440,n441,n442,n443,n444,n447,n448,n449,n450,n451,n453,n454,n455,n456,n457,n458,n459,n460,n461,n462,n463,n464,n465,n466,n467,n469,n470,n471,n472,n473,n474,n477,n478,n479,n480,n481,n483,n484,n485,n486,n487,n488,n489,n490,n491,n492,n493,n494,n495,n496,n497,n499,n500,n501,n502,n503,n504,n507,n508,n509,n510,n511,n513,n514,n515,n516,n517,n518,n519,n520,n521,n522,n523,n524,n525,n526,n527,n529,n530,n531,n532,n533,n534,n537,n538,n539,n540,n541,n543,n544,n545,n546,n547,n548,n549,n550,n551,n552,n553,n555,n556,n557,n558,n559,n560,n563,n564,n565,n566,n567,NS3,NS2,NS1,NS0,NS7,NS6,NS5,NS4,NS11,NS10,NS9,NS8,NS15,NS14,NS13,NS12,NS19,NS18,NS17,NS16,NS23,NS22,NS21,NS20,NS27,NS26,NS25,NS24,NS31,NS30,NS29,NS28;
not g0(n134,Clear);
not g1(n135,S3);
not g2(n136_1,S2);
not g3(n137,S1);
not g4(n138,S0);
not g5(n139,S7);
not g6(n140,S6);
not g7(n141_1,S5);
not g8(n142,S4);
not g9(n143,S11);
not g10(n144,S10);
not g11(n145,S9);
not g12(n146_1,S8);
not g13(n147,S15);
not g14(n148,S14);
not g15(n149,S13);
not g16(n150,S12);
not g17(n151_1,S19);
not g18(n152,S18);
not g19(n153,S17);
not g20(n154,S16);
not g21(n155,S23);
not g22(n156_1,S22);
not g23(n157,S21);
not g24(n158,S20);
not g25(n159,S27);
not g26(n160,S26);
not g27(n161_1,S25);
not g28(n162,S24);
not g29(n163,S31);
not g30(n164,S30);
not g31(n165,S29);
not g32(n166_1,S28);
and g33(n167,S29,S28);
not g34(n168,n167);
and g35(n169,S30,n167);
not g36(n170,n169);
and g37(W,S31,n169);
and g38(n172,X,n138);
and g39(n173,n137,n172);
and g40(n174,n136_1,n173);
and g41(n175,n135,n174);
and g42(n176_1,n142,n175);
and g43(n177,n141_1,n176_1);
and g44(n178,n140,n177);
and g45(n179,n139,n178);
and g46(n180,n146_1,n179);
and g47(n181_1,n145,n180);
and g48(n182,n144,n181_1);
and g49(n183,n143,n182);
and g50(n184,n150,n183);
and g51(n185,n149,n184);
and g52(n186_1,S14,n185);
and g53(n187,C_15,n186_1);
not g54(n188,n187);
and g55(n189,n148,n185);
and g56(n190,n147,n189);
and g57(n191_1,n154,n190);
and g58(n192,n153,n191_1);
and g59(n193,n152,n192);
and g60(n194,n151_1,n193);
and g61(n195,n158,n194);
and g62(n196_1,n157,n195);
and g63(n197,n156_1,n196_1);
and g64(n198,n155,n197);
and g65(n199,n162,n198);
and g66(n200,n161_1,n199);
and g67(n201_1,n160,n200);
and g68(n202,S27,n201_1);
and g69(n203,C_28,n202);
not g70(n204,n203);
and g71(n205,S10,n181_1);
and g72(n206_1,C_11,n205);
not g73(n207,n206_1);
and g74(n208,n204,n207);
and g75(n209,n188,n208);
and g76(n210,S9,n180);
and g77(n211_1,C_10,n210);
not g78(n212,n211_1);
and g79(n213,S2,n173);
and g80(n214,C_3,n213);
not g81(n215,n214);
and g82(n216_1,n212,n215);
and g83(n217,n209,n216_1);
and g84(n218,S16,n190);
and g85(n219,C_17,n218);
not g86(n220,n219);
and g87(n221_1,n159,n201_1);
and g88(n222,n166_1,n221_1);
and g89(n223,n165,n222);
and g90(n224,n164,n223);
and g91(n225,S31,n224);
and g92(n226_1,C_32,n225);
not g93(n227,n226_1);
and g94(n228,S23,n197);
and g95(n229,C_24,n228);
not g96(n230,n229);
and g97(n231_1,n227,n230);
and g98(n232,S22,n196_1);
and g99(n233,C_23,n232);
not g100(n234,n233);
and g101(n235,n231_1,n234);
and g102(n236,S13,n184);
and g103(n237,C_14,n236);
not g104(n238,n237);
and g105(n239,n235,n238);
and g106(n240,S25,n199);
and g107(n241,C_26,n240);
not g108(n242,n241);
and g109(n243,S1,n172);
and g110(n244,C_2,n243);
not g111(n245,n244);
and g112(n246,n242,n245);
and g113(n247,n239,n246);
and g114(n248,X,C_0);
not g115(n249,n248);
and g116(n250,S24,n198);
and g117(n251,C_25,n250);
not g118(n252,n251);
and g119(n253,n249,n252);
and g120(n254,S17,n191_1);
and g121(n255,C_18,n254);
not g122(n256,n255);
and g123(n257,S19,n193);
and g124(n258,C_20,n257);
not g125(n259,n258);
and g126(n260,n256,n259);
and g127(n261,S15,n189);
and g128(n262,C_16,n261);
not g129(n263,n262);
and g130(n264,S4,n175);
and g131(n265,C_5,n264);
not g132(n266,n265);
and g133(n267,n263,n266);
and g134(n268,n260,n267);
and g135(n269,n253,n268);
and g136(n270,n247,n269);
and g137(n271,n220,n270);
and g138(n272,S20,n194);
and g139(n273,C_21,n272);
not g140(n274,n273);
and g141(n275,S28,n221_1);
and g142(n276,C_29,n275);
not g143(n277,n276);
and g144(n278,S18,n192);
and g145(n279,C_19,n278);
not g146(n280,n279);
and g147(n281,n277,n280);
and g148(n282,S6,n177);
and g149(n283,C_7,n282);
not g150(n284,n283);
and g151(n285,n281,n284);
and g152(n286,S7,n178);
and g153(n287,C_8,n286);
not g154(n288,n287);
and g155(n289,S26,n200);
and g156(n290,C_27,n289);
not g157(n291,n290);
and g158(n292,n288,n291);
and g159(n293,n285,n292);
and g160(n294,S11,n182);
and g161(n295,C_12,n294);
not g162(n296,n295);
and g163(n297,S5,n176_1);
and g164(n298,C_6,n297);
not g165(n299,n298);
and g166(n300,n296,n299);
and g167(n301,n293,n300);
and g168(n302,n274,n301);
and g169(n303,S21,n195);
and g170(n304,C_22,n303);
not g171(n305,n304);
and g172(n306,X,S0);
and g173(n307,C_1,n306);
not g174(n308,n307);
and g175(n309,S29,n222);
and g176(n310,C_30,n309);
not g177(n311,n310);
and g178(n312,S30,n223);
and g179(n313,C_31,n312);
not g180(n314,n313);
and g181(n315,n311,n314);
and g182(n316,S3,n174);
and g183(n317,C_4,n316);
not g184(n318,n317);
and g185(n319,n315,n318);
and g186(n320,n308,n319);
and g187(n321,n305,n320);
and g188(n322,S12,n183);
and g189(n323,C_13,n322);
not g190(n324,n323);
and g191(n325,S8,n179);
and g192(n326,C_9,n325);
not g193(n327,n326);
and g194(n328,n324,n327);
and g195(n329,n321,n328);
and g196(n330,n302,n329);
and g197(n331,n271,n330);
and g198(n332,n217,n331);
not g199(Z,n332);
and g200(n334,X,n134);
and g201(n335,S0,n334);
and g202(n336,S1,n335);
and g203(n337,n135,S2);
and g204(n338,n336,n337);
not g205(n339,n338);
and g206(n340,S1,S0);
not g207(n341,n340);
and g208(n342,S2,n340);
not g209(n343,n342);
and g210(n344,n334,n343);
and g211(n345,S3,n344);
not g212(n346,n345);
and g213(n347,n339,n346);
not g214(NS3,n347);
and g215(n349,n334,n341);
and g216(n350,S2,n349);
not g217(n351,n350);
and g218(n352,n136_1,n336);
not g219(n353,n352);
and g220(n354,n351,n353);
not g221(NS2,n354);
and g222(NS0,n138,n334);
and g223(n357,S1,NS0);
not g224(n358,n357);
and g225(n359,n137,n335);
not g226(n360,n359);
and g227(n361,n358,n360);
not g228(NS1,n361);
and g229(n363,S3,n342);
and g230(n364,n134,n363);
and g231(n365,S4,n364);
and g232(n366,S5,n365);
and g233(n367,n139,S6);
and g234(n368,n366,n367);
not g235(n369,n368);
and g236(n370,S5,S4);
not g237(n371,n370);
and g238(n372,S6,n370);
not g239(n373,n372);
and g240(n374,n364,n373);
and g241(n375,S7,n374);
not g242(n376,n375);
and g243(n377,n369,n376);
not g244(NS7,n377);
and g245(n379,n364,n371);
and g246(n380,S6,n379);
not g247(n381,n380);
and g248(n382,n140,n366);
not g249(n383,n382);
and g250(n384,n381,n383);
not g251(NS6,n384);
and g252(NS4,n142,n364);
and g253(n387,S5,NS4);
not g254(n388,n387);
and g255(n389,n141_1,n365);
not g256(n390,n389);
and g257(n391,n388,n390);
not g258(NS5,n391);
and g259(n393,S7,n372);
and g260(n394,n134,n393);
and g261(n395,S8,n394);
and g262(n396,S9,n395);
and g263(n397,n143,S10);
and g264(n398,n396,n397);
not g265(n399,n398);
and g266(n400,S9,S8);
not g267(n401,n400);
and g268(n402,S10,n400);
not g269(n403,n402);
and g270(n404,n394,n403);
and g271(n405,S11,n404);
not g272(n406,n405);
and g273(n407,n399,n406);
not g274(NS11,n407);
and g275(n409,n394,n401);
and g276(n410,S10,n409);
not g277(n411,n410);
and g278(n412,n144,n396);
not g279(n413,n412);
and g280(n414,n411,n413);
not g281(NS10,n414);
and g282(NS8,n146_1,n394);
and g283(n417,S9,NS8);
not g284(n418,n417);
and g285(n419,n145,n395);
not g286(n420,n419);
and g287(n421,n418,n420);
not g288(NS9,n421);
and g289(n423,S11,n402);
and g290(n424,n134,n423);
and g291(n425,S12,n424);
and g292(n426,S13,n425);
and g293(n427,n147,S14);
and g294(n428,n426,n427);
not g295(n429,n428);
and g296(n430,S13,S12);
not g297(n431,n430);
and g298(n432,S14,n430);
not g299(n433,n432);
and g300(n434,n424,n433);
and g301(n435,S15,n434);
not g302(n436,n435);
and g303(n437,n429,n436);
not g304(NS15,n437);
and g305(n439,n424,n431);
and g306(n440,S14,n439);
not g307(n441,n440);
and g308(n442,n148,n426);
not g309(n443,n442);
and g310(n444,n441,n443);
not g311(NS14,n444);
and g312(NS12,n150,n424);
and g313(n447,S13,NS12);
not g314(n448,n447);
and g315(n449,n149,n425);
not g316(n450,n449);
and g317(n451,n448,n450);
not g318(NS13,n451);
and g319(n453,S15,n432);
and g320(n454,n134,n453);
and g321(n455,S16,n454);
and g322(n456,S17,n455);
and g323(n457,n151_1,S18);
and g324(n458,n456,n457);
not g325(n459,n458);
and g326(n460,S17,S16);
not g327(n461,n460);
and g328(n462,S18,n460);
not g329(n463,n462);
and g330(n464,n454,n463);
and g331(n465,S19,n464);
not g332(n466,n465);
and g333(n467,n459,n466);
not g334(NS19,n467);
and g335(n469,n454,n461);
and g336(n470,S18,n469);
not g337(n471,n470);
and g338(n472,n152,n456);
not g339(n473,n472);
and g340(n474,n471,n473);
not g341(NS18,n474);
and g342(NS16,n154,n454);
and g343(n477,S17,NS16);
not g344(n478,n477);
and g345(n479,n153,n455);
not g346(n480,n479);
and g347(n481,n478,n480);
not g348(NS17,n481);
and g349(n483,S19,n462);
and g350(n484,n134,n483);
and g351(n485,S20,n484);
and g352(n486,S21,n485);
and g353(n487,n155,S22);
and g354(n488,n486,n487);
not g355(n489,n488);
and g356(n490,S21,S20);
not g357(n491,n490);
and g358(n492,S22,n490);
not g359(n493,n492);
and g360(n494,n484,n493);
and g361(n495,S23,n494);
not g362(n496,n495);
and g363(n497,n489,n496);
not g364(NS23,n497);
and g365(n499,n484,n491);
and g366(n500,S22,n499);
not g367(n501,n500);
and g368(n502,n156_1,n486);
not g369(n503,n502);
and g370(n504,n501,n503);
not g371(NS22,n504);
and g372(NS20,n158,n484);
and g373(n507,S21,NS20);
not g374(n508,n507);
and g375(n509,n157,n485);
not g376(n510,n509);
and g377(n511,n508,n510);
not g378(NS21,n511);
and g379(n513,S23,n492);
and g380(n514,n134,n513);
and g381(n515,S24,n514);
and g382(n516,S25,n515);
and g383(n517,n159,S26);
and g384(n518,n516,n517);
not g385(n519,n518);
and g386(n520,S25,S24);
not g387(n521,n520);
and g388(n522,S26,n520);
not g389(n523,n522);
and g390(n524,n514,n523);
and g391(n525,S27,n524);
not g392(n526,n525);
and g393(n527,n519,n526);
not g394(NS27,n527);
and g395(n529,n514,n521);
and g396(n530,S26,n529);
not g397(n531,n530);
and g398(n532,n160,n516);
not g399(n533,n532);
and g400(n534,n531,n533);
not g401(NS26,n534);
and g402(NS24,n162,n514);
and g403(n537,S25,NS24);
not g404(n538,n537);
and g405(n539,n161_1,n515);
not g406(n540,n539);
and g407(n541,n538,n540);
not g408(NS25,n541);
and g409(n543,S27,n522);
and g410(n544,n134,n543);
and g411(n545,S28,n544);
and g412(n546,S29,n545);
and g413(n547,n163,S30);
and g414(n548,n546,n547);
not g415(n549,n548);
and g416(n550,n170,n544);
and g417(n551,S31,n550);
not g418(n552,n551);
and g419(n553,n549,n552);
not g420(NS31,n553);
and g421(n555,n168,n544);
and g422(n556,S30,n555);
not g423(n557,n556);
and g424(n558,n164,n546);
not g425(n559,n558);
and g426(n560,n557,n559);
not g427(NS30,n560);
and g428(NS28,n166_1,n544);
and g429(n563,S29,NS28);
not g430(n564,n563);
and g431(n565,n165,n545);
not g432(n566,n565);
and g433(n567,n564,n566);
not g434(NS29,n567);
always @(posedge clock) begin
S31<=NS31;
S30<=NS30;
S29<=NS29;
S28<=NS28;
S27<=NS27;
S26<=NS26;
S25<=NS25;
S24<=NS24;
S23<=NS23;
S22<=NS22;
S21<=NS21;
S20<=NS20;
S19<=NS19;
S18<=NS18;
S17<=NS17;
S16<=NS16;
S15<=NS15;
S14<=NS14;
S13<=NS13;
S12<=NS12;
S11<=NS11;
S10<=NS10;
S9<=NS9;
S8<=NS8;
S7<=NS7;
S6<=NS6;
S5<=NS5;
S4<=NS4;
S3<=NS3;
S2<=NS2;
S1<=NS1;
S0<=NS0;
end
endmodule
//State:00000000000000000000000010000000