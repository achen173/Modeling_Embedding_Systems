module ex3(clock,Rdy1RtHS1,Rdy2RtHS1,Rdy1BmHS1,Rdy2BmHS1,InDoneHS1,RtTSHS1,TpArrayHS1,OutputHS1,WantBmHS1,WantRtHS1,OutAvHS1,FullOHS1,FullIHS1,Prog_2,Prog_1,Prog_0,S26,S25,S22,S27,S14,S11,S17,S10,S13,S16,S6,S12,S19,S18,S15,S7,S9,S20,S28,S23,S8,S21,S24);
input clock;
input Rdy1RtHS1,Rdy2RtHS1,Rdy1BmHS1,Rdy2BmHS1,InDoneHS1,RtTSHS1,TpArrayHS1,OutputHS1,WantBmHS1,WantRtHS1,OutAvHS1,FullOHS1,FullIHS1,Prog_2,Prog_1,Prog_0;
output S26,S25,S22,S27,S14,S11,S17,S10,S13,S16,S6,S12,S19,S18,S15,S7,S9,S20,S28,S23,S8,S21,S24;
reg S0,S1,S2,S3,S4,S5,S6,S7,S8,S9,S10,S11,S12,S13,S14,S15,S16,S17,S18,S19,S20,S21,S22,S23,S24,S25,S26,S27,S28;
wire n127,n128,n129,n130_1,n131,n132,n133,n134_1,n135,n136,n137,n138_1,n139,n140,n141,n142_1,n143,n144,n145,n146_1,n147,n148,n149,n150_1,n151,n152,n153,n154_1,n155,n156,n157,n158_1,n159,n160,n161,n163,n164,n165,n166_1,n167,n168,n169,n170_1,n171,n173,n174_1,n175,n176,n177,n178_1,n179,n180,n181,n182_1,n183,n184,n185,n186_1,n187,n188,n189,n190_1,n191,n192,n193,n194_1,n195,n196,n197,n198_1,n199,n200,n201,n202,n203,n204,n205,n206,n207,n208,n209,n210,n211,n212,n213,n214,n215,n216,n217,n218,n219,n220,n221,n222,n223,n224,n225,n227,n228,n229,n230,n231,n232,n233,n234,n235,n236,n237,n238,n239,n240,n241,n242,n243,n244,n245,n246,n247,n248,n249,n250,n251,n252,n253,n254,n255,n256,n257,n258,n259,n260,n261,n262,n263,n264,n265,n266,n267,n268,n269,n270,n271,n272,n274,n275,n276,n277,n278,n279,n280,n281,n282,n283,n284,n285,n286,n287,n288,n289,n290,n291,n292,n293,n294,n295,n296,n297,n299,n300,n301,n302,n303,n304,n305,n306,n307,n308,n309,n310,n311,n312,n313,n314,n315,n316,n317,n318,n319,n320,n321,n322,n323,n324,n325,n326,n327,n328,n329,n331,n332,n333,n334,n335,n336,n337,n338,n339,n340,n341,n342,n343,n344,n345,n346,n347,n348,n349,n350,n351,n352,n353,n354,n355,n356,n357,n358,n359,n360,n361,n362,n363,n364,n365,n366,n367,n368,n369,n370,n371,n372,n373,n374,n375,n376,n377,n378,n379,n380,n381,n382,n383,n384,n385,n386,n387,n388,n389,n390,n391,n393,n394,n395,n396,n397,n398,n399,n400,n401,n402,n403,n404,n405,n406,n407,n408,n409,n410,n411,n412,n413,n414,n415,n416,n417,n418,n420,n421,n422,n423,n424,n425,n426,n427,n428,n429,n430,n431,n432,n433,n434,n435,n436,n438,n439,n440,n441,n442,n443,n444,n445,n446,n447,n448,n449,n450,n451,n452,n453,n454,n456,n457,n458,n459,n460,n461,n462,n463,n464,n465,n466,n467,n468,n469,n470,n471,n472,n473,n474,n475,n476,n477,n478,n479,n480,n481,n482,n484,n485,n486,n487,n488,n489,n490,n491,n492,n493,n494,n495,n496,n497,n498,n499,n500,n501,n502,n504,n506,n507,n508,n509,n510,n511,n512,n513,n514,n516,n517,n518,n519,n520,n521,n523,n524,n525,n526,n527,n528,n529,n530,n531,n532,n533,n534,n535,n536,n537,n539,n540,n541,n542,n543,n544,n545,n546,n547,n548,n549,n550,n552,n554,n555,n556,n557,n558,n559,n560,n561,n562,n563,n564,n565,n566,n567,n568,n569,n570,n571,n572,n573,n574,n576,n577,n578,n579,n580,n581,n582,n583,n584,n585,n586,n587,n588,n589,n590,n591,n592,n593,n594,n595,n596,n597,n599,n600,n601,n602,n603,n604,n605,n606,n607,n608,n609,n610,n611,n612,n613,n614,n615,n616,n617,n618,n619,n620,n621,n622,n623,n624,n626,n627,n628,n629,n630,n631,n632,n633,n634,n635,n636,n637,n638,n639,n640,n641,n642,n643,n644,n645,n646,n647,n648,n649,n652,n653,n654,n655,n656,n657,n658,n659,n660,n661,n662,n663,n664,n665,n667,n668,n669,n670,n671,n672,n673,n674,n678,n680,n681,n682,NS0,NS1,NS2,NS3,NS4,NS5,NS6,NS7,NS8,NS9,NS10,NS11,NS12,NS13,NS14,NS15,NS16,NS17,NS18,NS19,NS20,NS21,NS22,NS23,NS24,NS25,NS26,NS27,NS28;
not g0(n127,Rdy1RtHS1);
not g1(n128,Rdy2RtHS1);
not g2(n129,Rdy1BmHS1);
not g3(n130_1,Rdy2BmHS1);
not g4(n131,InDoneHS1);
not g5(n132,TpArrayHS1);
not g6(n133,WantBmHS1);
not g7(n134_1,WantRtHS1);
not g8(n135,OutAvHS1);
not g9(n136,FullOHS1);
not g10(n137,FullIHS1);
not g11(n138_1,Prog_2);
not g12(n139,Prog_1);
not g13(n140,Prog_0);
not g14(n141,S0);
not g15(n142_1,S1);
not g16(n143,S2);
not g17(n144,S3);
not g18(n145,S4);
not g19(n146_1,S5);
and g20(n147,S0,n143);
and g21(n148,n144,n147);
and g22(n149,n136,n137);
not g23(n150_1,n149);
and g24(n151,n142_1,n150_1);
and g25(n152,n148,n151);
and g26(n153,S5,n152);
not g27(n154_1,n153);
and g28(n155,n142_1,n148);
and g29(n156,n129,n155);
and g30(n157,n127,n156);
not g31(n158_1,n157);
and g32(n159,n154_1,n158_1);
and g33(n160,n145,n148);
and g34(n161,S1,n146_1);
and g35(NS14,n160,n161);
not g36(n163,NS14);
and g37(n164,n138_1,n139);
not g38(n165,n164);
and g39(n166_1,RtTSHS1,n143);
not g40(n167,n166_1);
and g41(n168,n141,n142_1);
and g42(n169,S3,n146_1);
and g43(n170_1,n168,n169);
and g44(n171,n145,n170_1);
and g45(NS11,n166_1,n171);
and g46(n173,n165,NS11);
not g47(n174_1,n173);
and g48(n175,n163,n174_1);
and g49(n176,n159,n175);
and g50(n177,n145,n146_1);
not g51(n178_1,n177);
and g52(n179,S4,S5);
not g53(n180,n179);
and g54(n181,n178_1,n180);
and g55(n182_1,S3,n147);
and g56(n183,n181,n182_1);
not g57(n184,n183);
and g58(n185,Prog_2,n160);
not g59(n186_1,n185);
and g60(n187,n146_1,n185);
not g61(n188,n187);
and g62(n189,n184,n188);
and g63(n190_1,Rdy1BmHS1,Rdy2BmHS1);
not g64(n191,n190_1);
and g65(n192,n140,n160);
not g66(n193,n192);
and g67(n194_1,n145,S5);
and g68(n195,n147,n194_1);
not g69(n196,n195);
and g70(n197,n193,n196);
not g71(n198_1,n197);
and g72(n199,n191,n198_1);
not g73(n200,n199);
and g74(n201,Prog_2,n152);
not g75(n202,n201);
and g76(n203,n200,n202);
and g77(n204,n138_1,n142_1);
not g78(n205,n204);
and g79(n206,n181,n204);
and g80(n207,n147,n206);
not g81(n208,n207);
and g82(n209,Rdy1RtHS1,Rdy2RtHS1);
not g83(n210,n209);
and g84(n211,n146_1,n148);
and g85(n212,Prog_0,n211);
not g86(n213,n212);
and g87(n214,S4,n146_1);
and g88(n215,n143,n214);
and g89(n216,S0,n215);
not g90(n217,n216);
and g91(n218,n213,n217);
not g92(n219,n218);
and g93(n220,n210,n219);
not g94(n221,n220);
and g95(n222,n208,n221);
and g96(n223,n203,n222);
and g97(n224,n189,n223);
and g98(n225,n176,n224);
not g99(NS0,n225);
and g100(n227,n128,n214);
not g101(n228,n227);
and g102(n229,n130_1,n194_1);
not g103(n230,n229);
and g104(n231,n228,n230);
not g105(n232,n231);
and g106(n233,n147,n232);
not g107(n234,n233);
and g108(n235,n184,n234);
not g109(n236,n235);
and g110(n237,S1,n236);
not g111(n238,n237);
and g112(n239,Rdy1BmHS1,n130_1);
not g113(n240,n239);
and g114(n241,WantBmHS1,n240);
not g115(n242,n241);
and g116(n243,n142_1,n149);
and g117(n244,n185,n243);
and g118(n245,n146_1,n244);
and g119(n246,Rdy2RtHS1,n245);
not g120(n247,n246);
and g121(n248,n242,n246);
and g122(n249,Prog_0,n248);
not g123(n250,n249);
and g124(n251,n238,n250);
and g125(n252,n131,NS14);
not g126(n253,n252);
and g127(n254,Rdy1RtHS1,n128);
not g128(n255,n254);
and g129(n256,WantRtHS1,n255);
not g130(n257,n256);
and g131(n258,n245,n257);
and g132(n259,n139,n140);
not g133(n260,n259);
and g134(n261,Prog_1,Prog_0);
not g135(n262,n261);
and g136(n263,n260,n262);
not g137(n264,n263);
and g138(n265,Rdy2BmHS1,n263);
not g139(n266,n265);
and g140(n267,n241,n266);
not g141(n268,n267);
and g142(n269,n258,n268);
not g143(n270,n269);
and g144(n271,n253,n270);
and g145(n272,n251,n271);
not g146(NS1,n272);
and g147(n274,n146_1,n149);
and g148(n275,n190_1,n274);
not g149(n276,n275);
and g150(n277,n143,n276);
not g151(n278,n277);
and g152(n279,n145,n278);
and g153(n280,n168,n279);
and g154(n281,n144,n280);
not g155(n282,n281);
and g156(n283,S2,n168);
and g157(n284,n194_1,n283);
not g158(n285,n284);
and g159(n286,n144,n283);
and g160(n287,S5,n286);
not g161(n288,n287);
and g162(n289,n132,n287);
not g163(n290,n289);
and g164(n291,n285,n290);
and g165(n292,S4,n170_1);
not g166(n293,n292);
and g167(n294,S2,n292);
not g168(n295,n294);
and g169(n296,n291,n295);
and g170(n297,n282,n296);
not g171(NS2,n297);
and g172(n299,n136,Prog_2);
and g173(n300,n137,n299);
not g174(n301,n300);
and g175(n302,n142_1,n301);
not g176(n303,n302);
and g177(n304,S4,n303);
and g178(n305,n211,n304);
and g179(n306,n254,n305);
not g180(n307,n306);
and g181(n308,S5,n303);
and g182(n309,n160,n308);
and g183(n310,n239,n309);
not g184(n311,n310);
and g185(n312,n307,n311);
and g186(n313,n142_1,n145);
and g187(n314,n143,n144);
and g188(n315,n313,n314);
and g189(n316,n141,n275);
and g190(n317,n315,n316);
not g191(n318,n317);
and g192(n319,n170_1,n167);
not g193(n320,n319);
and g194(n321,n318,n320);
and g195(n322,S4,n287);
not g196(n323,n322);
and g197(n324,n131,n183);
not g198(n325,n324);
and g199(n326,n323,n325);
and g200(n327,n321,n326);
and g201(n328,n312,n327);
and g202(n329,n293,n328);
not g203(NS3,n329);
and g204(n331,Rdy2BmHS1,WantBmHS1);
and g205(n332,Prog_2,n211);
not g206(n333,n332);
and g207(n334,Rdy1RtHS1,n332);
and g208(n335,n243,n334);
and g209(n336,n145,n335);
not g210(n337,n336);
and g211(n338,n247,n337);
not g212(n339,n338);
and g213(n340,n331,n339);
not g214(n341,n340);
and g215(n342,n134_1,n245);
not g216(n343,n342);
and g217(n344,n331,n342);
not g218(n345,n344);
and g219(n346,n341,n345);
and g220(n347,n131,n138_1);
not g221(n348,n347);
and g222(n349,Prog_2,n150_1);
not g223(n350,n349);
and g224(n351,n348,n350);
not g225(n352,n351);
and g226(n353,n142_1,n352);
not g227(n354,n353);
and g228(n355,n144,n354);
and g229(n356,n205,n210);
not g230(n357,n356);
and g231(n358,n355,n357);
not g232(n359,n358);
and g233(n360,n216,n359);
not g234(n361,n360);
and g235(n362,n129,Rdy2BmHS1);
and g236(n363,n309,n362);
not g237(n364,n363);
and g238(n365,n361,n364);
and g239(n366,n346,n365);
and g240(n367,n140,n239);
not g241(n368,n367);
and g242(n369,Prog_0,n254);
not g243(n370,n369);
and g244(n371,n368,n370);
not g245(n372,n371);
and g246(n373,n138_1,n211);
and g247(n374,n137,n373);
and g248(n375,FullOHS1,n374);
and g249(n376,n313,n375);
and g250(n377,n372,n376);
not g251(n378,n377);
and g252(n379,n131,n294);
not g253(n380,n379);
and g254(n381,n378,n380);
and g255(n382,S4,n153);
not g256(n383,n382);
and g257(n384,n142_1,n215);
and g258(n385,S3,n384);
and g259(n386,n210,n385);
not g260(n387,n386);
and g261(n388,n383,n387);
and g262(n389,n381,n388);
and g263(n390,n288,n389);
and g264(n391,n366,n390);
not g265(NS4,n391);
and g266(n393,n129,n130_1);
not g267(n394,n393);
and g268(n395,WantBmHS1,n393);
not g269(n396,n395);
and g270(n397,WantRtHS1,n246);
and g271(n398,n396,n397);
not g272(n399,n398);
and g273(n400,n383,n399);
and g274(n401,n313,n373);
not g275(n402,n401);
and g276(n403,n136,n401);
and g277(n404,n372,n403);
not g278(n405,n404);
and g279(n406,n282,n405);
and g280(n407,n127,Rdy2RtHS1);
and g281(n408,n305,n407);
not g282(n409,n408);
and g283(n410,n191,n205);
not g284(n411,n410);
and g285(n412,n355,n411);
not g286(n413,n412);
and g287(n414,n195,n413);
not g288(n415,n414);
and g289(n416,n409,n415);
and g290(n417,n406,n416);
and g291(n418,n400,n417);
not g292(NS5,n418);
and g293(n420,n182_1,n214);
not g294(n421,n420);
and g295(n422,n163,n421);
and g296(n423,n138_1,n194_1);
not g297(n424,n423);
and g298(n425,n142_1,n147);
and g299(n426,n423,n425);
not g300(n427,n426);
and g301(n428,Prog_0,n144);
and g302(n429,n426,n428);
not g303(n430,n429);
and g304(n431,n138_1,S0);
and g305(n432,n384,n431);
and g306(n433,Prog_0,n432);
not g307(n434,n433);
and g308(n435,n430,n434);
and g309(n436,n422,n435);
not g310(NS6,n436);
and g311(n438,n182_1,n194_1);
not g312(n439,n438);
and g313(n440,n163,n439);
and g314(n441,n144,n432);
not g315(n442,n441);
and g316(n443,n427,n442);
not g317(n444,n443);
and g318(n445,n140,n444);
not g319(n446,n445);
and g320(n447,n144,S4);
not g321(n448,n447);
and g322(n449,n146_1,n448);
and g323(n450,n283,n449);
not g324(n451,n450);
and g325(n452,n446,n451);
and g326(n453,n288,n452);
and g327(n454,n440,n453);
not g328(NS7,n454);
and g329(n456,n128,n335);
not g330(n457,n456);
and g331(n458,n242,n456);
and g332(n459,WantRtHS1,n458);
not g333(n460,n459);
and g334(n461,n307,n460);
and g335(n462,n127,n128);
not g336(n463,n462);
and g337(n464,n210,n463);
and g338(n465,n401,n464);
and g339(n466,FullOHS1,FullIHS1);
not g340(n467,n466);
and g341(n468,Prog_0,n467);
and g342(n469,n465,n468);
not g343(n470,n469);
and g344(n471,n127,n136);
and g345(n472,n137,n155);
and g346(n473,n129,n472);
and g347(n474,n179,n473);
and g348(n475,n471,n474);
not g349(n476,n475);
and g350(n477,n470,n476);
and g351(n478,n461,n477);
and g352(n479,n209,n292);
and g353(n480,n143,n479);
not g354(n481,n480);
and g355(n482,n478,n481);
not g356(NS8,n482);
and g357(n484,n146_1,n204);
and g358(n485,n192,n484);
and g359(n486,n239,n485);
not g360(n487,n486);
and g361(n488,n362,n485);
not g362(n489,n488);
and g363(n490,n487,n489);
not g364(n491,n490);
and g365(n492,n467,n491);
not g366(n493,n492);
and g367(n494,n476,n493);
and g368(n495,n244,n257);
and g369(n496,n239,n495);
not g370(n497,n496);
and g371(n498,WantBmHS1,n496);
not g372(n499,n498);
and g373(n500,n318,n499);
and g374(n501,n311,n500);
and g375(n502,n494,n501);
not g376(NS9,n502);
and g377(n504,n288,n451);
not g378(NS10,n504);
and g379(n506,S0,n385);
not g380(n507,n506);
and g381(n508,Prog_0,NS14);
not g382(n509,n508);
and g383(n510,n507,n509);
and g384(n511,n140,n432);
not g385(n512,n511);
and g386(n513,n430,n512);
and g387(n514,n510,n513);
not g388(NS12,n514);
and g389(n516,Prog_1,NS14);
not g390(n517,n516);
and g391(n518,n142_1,n183);
not g392(n519,n518);
and g393(n520,n208,n519);
and g394(n521,n517,n520);
not g395(NS13,n521);
and g396(n523,Prog_2,NS11);
not g397(n524,n523);
and g398(n525,n318,n524);
and g399(n526,Rdy1RtHS1,n227);
not g400(n527,n526);
and g401(n528,Rdy1BmHS1,n229);
not g402(n529,n528);
and g403(n530,n527,n529);
not g404(n531,n530);
and g405(n532,n472,n531);
and g406(n533,n299,n532);
not g407(n534,n533);
and g408(n535,n402,n476);
and g409(n536,n534,n535);
and g410(n537,n525,n536);
not g411(NS15,n537);
and g412(n539,S3,n181);
not g413(n540,n539);
and g414(n541,n424,n540);
not g415(n542,n541);
and g416(n543,n425,n542);
not g417(n544,n543);
and g418(n545,n295,n544);
and g419(n546,n145,n286);
not g420(n547,n546);
and g421(n548,n163,n547);
and g422(n549,n288,n548);
and g423(n550,n545,n549);
not g424(NS16,n550);
and g425(n552,n163,n442);
not g426(NS17,n552);
and g427(n554,Prog_2,n315);
and g428(n555,n146_1,n554);
not g429(n556,n555);
and g430(n557,n192,n467);
not g431(n558,n557);
and g432(n559,n186_1,n558);
not g433(n560,n559);
and g434(n561,n130_1,n560);
not g435(n562,n561);
and g436(n563,n556,n562);
and g437(n564,n212,n467);
not g438(n565,n564);
and g439(n566,n333,n565);
not g440(n567,n566);
and g441(n568,n128,n567);
not g442(n569,n568);
and g443(n570,n177,n168);
not g444(n571,n570);
and g445(n572,n569,n571);
and g446(n573,n288,n572);
and g447(n574,n563,n573);
not g448(NS18,n574);
and g449(n576,n140,n373);
and g450(n577,Rdy2BmHS1,n136);
and g451(n578,n576,n577);
not g452(n579,n578);
and g453(n580,S5,n156);
not g454(n581,n580);
and g455(n582,n579,n581);
and g456(n583,Rdy2RtHS1,Prog_0);
not g457(n584,n583);
and g458(n585,n129,n140);
not g459(n586,n585);
and g460(n587,n584,n586);
not g461(n588,n587);
and g462(n589,n374,n588);
not g463(n590,n589);
and g464(n591,n571,n590);
and g465(n592,n212,n471);
and g466(n593,n138_1,n592);
not g467(n594,n593);
and g468(n595,n288,n594);
and g469(n596,n591,n595);
and g470(n597,n582,n596);
not g471(NS19,n597);
and g472(n599,S3,n177);
not g473(n600,n599);
and g474(n601,n144,n179);
and g475(n602,TpArrayHS1,n601);
not g476(n603,n602);
and g477(n604,n600,n603);
not g478(n605,n604);
and g479(n606,n283,n605);
not g480(n607,n606);
and g481(n608,n343,n457);
not g482(n609,n608);
and g483(n610,n133,n609);
not g484(n611,n610);
and g485(n612,n497,n611);
and g486(n613,Prog_0,n403);
and g487(n614,n464,n613);
not g488(n615,n614);
and g489(n616,n191,n394);
and g490(n617,n485,n616);
and g491(n618,n136,n617);
not g492(n619,n618);
and g493(n620,n615,n619);
and g494(n621,n476,n534);
and g495(n622,n620,n621);
and g496(n623,n612,n622);
and g497(n624,n607,n623);
not g498(NS20,n624);
and g499(n626,n138_1,Prog_0);
and g500(n627,n127,FullOHS1);
and g501(n628,n626,n627);
not g502(n629,n628);
and g503(n630,n133,n140);
and g504(n631,n299,n630);
and g505(n632,WantRtHS1,n631);
not g506(n633,n632);
and g507(n634,n629,n633);
not g508(n635,n634);
and g509(n636,Rdy2RtHS1,n635);
and g510(n637,n472,n636);
and g511(n638,n177,n637);
not g512(n639,n638);
and g513(n640,n264,n344);
not g514(n641,n640);
and g515(n642,n639,n641);
and g516(n643,n140,n616);
not g517(n644,n643);
and g518(n645,n370,n644);
not g519(n646,n645);
and g520(n647,n376,n646);
not g521(n648,n647);
and g522(n649,n642,n648);
not g523(NS21,n649);
and g524(NS22,n135,n150_1);
and g525(n652,n136,n488);
not g526(n653,n652);
and g527(n654,n407,n613);
not g528(n655,n654);
and g529(n656,n476,n655);
and g530(n657,OutputHS1,NS14);
not g531(n658,n657);
and g532(n659,n544,n658);
not g533(n660,n659);
and g534(n661,InDoneHS1,n660);
not g535(n662,n661);
and g536(n663,n607,n662);
and g537(n664,n656,n663);
and g538(n665,n653,n664);
not g539(NS23,n665);
and g540(n667,InDoneHS1,n441);
not g541(n668,n667);
and g542(n669,n639,n668);
and g543(n670,n137,n488);
and g544(n671,FullOHS1,n670);
not g545(n672,n671);
and g546(n673,n641,n672);
and g547(n674,n669,n673);
not g548(NS24,n674);
and g549(NS25,n135,FullIHS1);
and g550(NS26,n135,n137);
and g551(n678,S2,n144);
and g552(NS27,n570,n678);
and g553(n680,n397,n630);
not g554(n681,n680);
and g555(n682,n641,n681);
not g556(NS28,n682);
always @ (posedge clock) begin
S28<=NS28;
S27<=NS27;
S26<=NS26;
S25<=NS25;
S24<=NS24;
S23<=NS23;
S22<=NS22;
S21<=NS21;
S20<=NS20;
S19<=NS19;
S18<=NS18;
S17<=NS17;
S16<=NS16;
S15<=NS15;
S14<=NS14;
S13<=NS13;
S12<=NS12;
S11<=NS11;
S10<=NS10;
S9<=NS9;
S8<=NS8;
S7<=NS7;
S6<=NS6;
S5<=NS5;
S4<=NS4;
S3<=NS3;
S2<=NS2;
S1<=NS1;
S0<=NS0;
end
endmodule
//State:00000000010110110000011000001